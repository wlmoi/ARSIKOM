// Praktikum EL3011 Arsitektur Sistem Komputer
// Modul      : 2
// Percobaan  : 1
// Tanggal    : 19 November 2025
// Nama (NIM) 1 : William Anthony (13223048)
// Nama (NIM) 2 : Agita Trinanda Ilmi (13223003)
// Nama File  : mux2to1_rv32i.v
// Deskripsi  : Desain multiplexer 2-ke-1 generik 32-bit

module mux2to1_rv32i #(parameter WIDTH = 32) (
    input  wire [WIDTH-1:0] in0, // Input pertama
    input  wire [WIDTH-1:0] in1, // Input kedua
    input  wire sel,             // Sinyal seleksi (0 = in0, 1 = in1)
    output wire [WIDTH-1:0] out  // Output yang dipilih
);
    assign out = sel ? in1 : in0; // Logika multiplexer
endmodule
